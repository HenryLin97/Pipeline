library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
--ע����ͳһ�� 0 ��ʾʹ��
--��1��ʾ��ʹ��
entity NewMemoryTest is
	Port( clk : in std_logic;
			rst : in std_logic;
			keep_im : in std_logic; --when this is 1, keep imOut!
			--DM
			dmControl : in std_logic_vector(2 downto 0);-- 001 �� 010 д
			--dmWrite: in std_logic; --��0��ʾ��Ҫд���Ӧ��ram
			--dmRead : in std_logic; --��0��ʾ��Ҫ��ȡ��Ӧ��ram
			dmAddr : in std_logic_vector(15 downto 0); --����ram�õĵ�ַ��ע����������õ������ַ
			dmIn : in std_logic_vector(15 downto 0);		--д�ڴ�ʱ��Ҫд��ram1������
			dmOut : out std_logic_vector(15 downto 0);	--��DMʱ��������������/�����Ĵ���״̬
			--IM
			--WriteIM : in std_logic;
			--imRead : in std_logic;
			imAddr : in std_logic_vector(15 downto 0);
			--imIn:	in std_logic_vector(15 downto 0);
			imOut:	out std_logic_vector(15 downto 0);
			Memory_PCOut : out std_logic_vector(15 downto 0);
			--UART�����ź�  
			ram1_oe, ram1_we, ram1_en : out STD_LOGIC;
			ram2_oe, ram2_we, ram2_en : out STD_LOGIC;
			ram1_addr, ram2_addr : out STD_LOGIC_VECTOR(17 downto 0); --����ram�ĵ�ַ����
			ram1_data, ram2_data : inout STD_LOGIC_VECTOR(15 downto 0); --����ram����������
			data_ready : in std_logic;
			tbre : in std_logic;
			tsre : in std_logic;
			wrn : out std_logic;
			rdn : out std_logic;
			--�����ź�
			display_im : out std_logic_vector(15 downto 0);
			display_dm : out std_logic_vector(15 downto 0);
			--��������ź�
--			dm_data_ready : out std_logic;
--			im_data_ready : out std_logic;
			stall_im : in std_logic;
			stall_dm : in std_logic;
			flush : in std_logic;
			--�������
			req_stall_im :out std_logic;
			req_stall_dm :out std_logic
			);
end NewMemoryTest;

architecture Behavioral of NewMemoryTest is
shared variable count: INTEGER range 0 to 10 := 0;
Constant border_position : integer range 0 to 65536:=32768;--0x8000
Constant chuankou_position : integer range 0 to 65536:=48896;--0xBF00
Constant chuankou_status_position : integer range 0 to 65536:=48897; --0xBF01
shared variable position : integer range 0 to 65536:=0;
type dm_target_type is (RAM1,RAM2,CHUANKOU,CHUANKOU_STATUS);
shared variable dm_target : dm_target_type;
signal im_state : std_logic := '0'; --use to simulate memory stop
signal dm_state : std_logic := '0'; --use to simulate memory stop
signal current_data : std_logic_vector(15 downto 0):=(others => '0');
shared variable dmout_temp : std_logic_vector(15 downto 0);
shared variable imout_temp : std_logic_vector(15 downto 0);
--
shared variable state_keep : std_logic :='0';
shared variable dmcontrol_state : std_logic_vector(2 downto 0);
shared variable keep_im_state : std_logic ;
begin
	process(clk, rst)
	begin
		if(rst = '0') then
			ram1_oe <= '1';
			ram1_we <= '1';
			ram1_en <= '1';
			ram2_oe <= '1';
			ram2_we <= '1';
			ram2_en <= '1';
			wrn <= '1';
			rdn <= '1';
			--req_stall_im <= '0';
			req_stall_dm <= '0';
			--dm_data_ready <= '1';
			--im_data_ready <= '1';
			imOut_temp := "0000100000000000";
			dmOut_temp := "1111111111111111";
			Memory_PCOut <= (others=>'1');
		elsif(rising_edge(clk)) then
			--imOut <= "0100000101000001"; -- instruction
			--get dm postion 
			if(state_keep = '0') then
				position := CONV_INTEGER(dmAddr);
				if(position < border_position) then
					dm_target:= RAM2; --IM
				elsif(position = chuankou_position) then
					dm_target:= CHUANKOU;
				elsif(position = chuankou_status_position) then
					dm_target:= CHUANKOU_STATUS;
				else
					dm_target:= RAM1; --DM
				end if;
				dmControl_state := dmcontrol;
				keep_im_state := keep_im;
			else
				state_keep := '0';
			end if;
			Memory_PCOut <= imAddr;
			if(dmControl_state = "001")then	--read
				case dm_target is
					when RAM1 =>
						dmOut_temp := "0010000000000001";
					when RAM2 =>
						dmOut_temp := "0010000000000010";
					when CHUANKOU =>--BF00
						dmOut_temp := "0000000001010010";
						state_keep := '1';
					when CHUANKOU_STATUS =>
						--dmOut_temp := "0010000000000100";
						dmOut_temp := "0100000000000101";
				end case;
				 --memory value
			elsif(dmControl_state = "010")then  --write
				case dm_target is
					when RAM1 =>
						dmOut_temp := "0100000000000001";
					when RAM2 =>
						dmOut_temp := "0100000000000010";
					when CHUANKOU =>--BF00
						dmOut_temp := "0100000000000011";
						state_keep := '1';
						--req_stall_dm <= '1';
					when CHUANKOU_STATUS =>
						dmOut_temp := "0100000000000100";
						--dmOut_temp := "0100000000000101";
				end case;
			else
			end if;
			if (keep_im_state = '0') then
				if (im_state = '1') then
					imOut_temp := "0100001000100001";
					--req_stall_im <= '0';
					im_state <= '0';
				else
				case imAddr is
--				when "0000000000000000"=>
--    imOut_temp :="0000000000000000";
when "0000000000000000"=>
	imOut_temp := "0110100000000001";
when "0000000000000001"=>
    imOut_temp :="0110100100000001";
when "0000000000000010"=>
    imOut_temp :="1110100000101010";
when "0000000000000011"=>
    imOut_temp :="0110000000110010";
--when "0000000000000001"=>
--    imOut_temp :="0000000000000000";
--when "0000000000000010"=>
--    imOut_temp :="0000100000000000";
--when "0000000000000011"=>
--    imOut_temp :="0001000001100001";
when "0000000000000100"=>
    imOut_temp :="0000100000000000";
when "0000000000000101"=>
    imOut_temp :="0000100000000000";
when "0000000000000110"=>
    imOut_temp :="0000100000000000";
when "0000000000000111"=>
    imOut_temp :="0000100000000000";
when "0000000000001000"=>
    imOut_temp :="0110111010111111";
when "0000000000001001"=>
    imOut_temp :="0011011011000000";
when "0000000000001010"=>
    imOut_temp :="0100111000010000";
when "0000000000001011"=>
    imOut_temp :="1101111000000000";
when "0000000000001100"=>
    imOut_temp :="1101111000100001";
when "0000000000001101"=>
    imOut_temp :="1101111001000010";
when "0000000000001110"=>
    imOut_temp :="1101111010000100";
when "0000000000001111"=>
    imOut_temp :="1101111010100101";
when "0000000000010000"=>
    imOut_temp :="1001000100000000";
when "0000000000010001"=>
    imOut_temp :="0110001100000001";
when "0000000000010010"=>
    imOut_temp :="0110100011111111";
when "0000000000010011"=>
    imOut_temp :="1110100100001100";
when "0000000000010100"=>
    imOut_temp :="1001001000000000";
when "0000000000010101"=>
    imOut_temp :="0110001100000001";
when "0000000000010110"=>
    imOut_temp :="0110001111111111";
when "0000000000010111"=>
    imOut_temp :="1101001100000000";
when "0000000000011000"=>
    imOut_temp :="0110001111111111";
when "0000000000011001"=>
    imOut_temp :="1101011100000000";
when "0000000000011010"=>
    imOut_temp :="0110101100001111";
when "0000000000011011"=>
    imOut_temp :="1110111101000000";
when "0000000000011100"=>
    imOut_temp :="0100111100000011";
when "0000000000011101"=>
    imOut_temp :="0000100000000000";
when "0000000000011110"=>
    imOut_temp :="0001000010101100";
when "0000000000011111"=>
    imOut_temp :="0000100000000000";
when "0000000000100000"=>
    imOut_temp :="0110111010111111";
when "0000000000100001"=>
    imOut_temp :="0011011011000000";
when "0000000000100010"=>
    imOut_temp :="1101111001100000";
when "0000000000100011"=>
    imOut_temp :="0000100000000000";
when "0000000000100100"=>
    imOut_temp :="0110111010111111";
when "0000000000100101"=>
    imOut_temp :="0011011011000000";
when "0000000000100110"=>
    imOut_temp :="0100111000010000";
when "0000000000100111"=>
    imOut_temp :="0110100000000000";
when "0000000000101000"=>
    imOut_temp :="1110100000101010";
when "0000000000101001"=>
    imOut_temp :="0110000100000010";
when "0000000000101010"=>
    imOut_temp :="0000100000000000";
when "0000000000101011"=>
    imOut_temp :="1001111010000111";
when "0000000000101100"=>
    imOut_temp :="0110100000100000";
when "0000000000101101"=>
    imOut_temp :="1110100000101010";
when "0000000000101110"=>
    imOut_temp :="0110000100000010";
when "0000000000101111"=>
    imOut_temp :="0000100000000000";
when "0000000000110000"=>
    imOut_temp :="1001111010001000";
when "0000000000110001"=>
    imOut_temp :="0110100000010000";
when "0000000000110010"=>
    imOut_temp :="1110100000101010";
when "0000000000110011"=>
    imOut_temp :="0110000100000010";
when "0000000000110100"=>
    imOut_temp :="0000100000000000";
when "0000000000110101"=>
    imOut_temp :="1001111010001001";
when "0000000000110110"=>
    imOut_temp :="0000100000000000";
when "0000000000110111"=>
    imOut_temp :="1001111010100110";
when "0000000000111000"=>
    imOut_temp :="1110110010100010";
when "0000000000111001"=>
    imOut_temp :="0110000100001011";
when "0000000000111010"=>
    imOut_temp :="0000100000000000";
when "0000000000111011"=>
    imOut_temp :="1101111010000110";
when "0000000000111100"=>
    imOut_temp :="1110111101000000";
when "0000000000111101"=>
    imOut_temp :="0100111100000011";
when "0000000000111110"=>
    imOut_temp :="0000100000000000";
when "0000000000111111"=>
    imOut_temp :="0001000010001011";
when "0000000001000000"=>
    imOut_temp :="0000100000000000";
when "0000000001000001"=>
    imOut_temp :="0110111010111111";
when "0000000001000010"=>
    imOut_temp :="0011011011000000";
when "0000000001000011"=>
    imOut_temp :="1101111000100000";
when "0000000001000100"=>
    imOut_temp :="0000100000000000";
when "0000000001000101"=>
    imOut_temp :="0000100000000000";
when "0000000001000110"=>
    imOut_temp :="0110101100001111";
when "0000000001000111"=>
    imOut_temp :="1110111101000000";
when "0000000001001000"=>
    imOut_temp :="0100111100000011";
when "0000000001001001"=>
    imOut_temp :="0000100000000000";
when "0000000001001010"=>
    imOut_temp :="0001000010000000";
when "0000000001001011"=>
    imOut_temp :="0000100000000000";
when "0000000001001100"=>
    imOut_temp :="0110111010111111";
when "0000000001001101"=>
    imOut_temp :="0011011011000000";
when "0000000001001110"=>
    imOut_temp :="1101111001100000";
when "0000000001001111"=>
    imOut_temp :="0000100000000000";
when "0000000001010000"=>
    imOut_temp :="0100001011000000";
when "0000000001010001"=>
    imOut_temp :="1111001100000000";
when "0000000001010010"=>
    imOut_temp :="0110100010000000";
when "0000000001010011"=>
    imOut_temp :="0011000000000000";
when "0000000001010100"=>
    imOut_temp :="1110101100001101";
when "0000000001010101"=>
    imOut_temp :="0110111110111111";
when "0000000001010110"=>
    imOut_temp :="0011011111100000";
when "0000000001010111"=>
    imOut_temp :="0100111100010000";
when "0000000001011000"=>
    imOut_temp :="1001111100000000";
when "0000000001011001"=>
    imOut_temp :="1001111100100001";
when "0000000001011010"=>
    imOut_temp :="1001111101000010";
when "0000000001011011"=>
    imOut_temp :="1001111110000100";
when "0000000001011100"=>
    imOut_temp :="1001111110100101";
when "0000000001011101"=>
    imOut_temp :="1001011100000000";
when "0000000001011110"=>
    imOut_temp :="0110001100000001";
when "0000000001011111"=>
    imOut_temp :="0110001100000001";
when "0000000001100000"=>
    imOut_temp :="0000100000000000";
when "0000000001100001"=>
    imOut_temp :="1111001100000001";
when "0000000001100010"=>
    imOut_temp :="1110111000000000";
when "0000000001100011"=>
    imOut_temp :="1001001111111111";
when "0000000001100100"=>
    imOut_temp :="0000100000000000";
when "0000000001100101"=>
    imOut_temp :="0110100000000111";
when "0000000001100110"=>
    imOut_temp :="1111000000000001";
when "0000000001100111"=>
    imOut_temp :="0110100010111111";
when "0000000001101000"=>
    imOut_temp :="0011000000000000";
when "0000000001101001"=>
    imOut_temp :="0100100000010000";
when "0000000001101010"=>
    imOut_temp :="0110010000000000";
when "0000000001101011"=>
    imOut_temp :="0000100000000000";
when "0000000001101100"=>
    imOut_temp :="0110111010111111";
when "0000000001101101"=>
    imOut_temp :="0011011011000000";
when "0000000001101110"=>
    imOut_temp :="0100111000010000";
when "0000000001101111"=>
    imOut_temp :="0110100000000000";
when "0000000001110000"=>
    imOut_temp :="1101111000000000";
when "0000000001110001"=>
    imOut_temp :="1101111000000001";
when "0000000001110010"=>
    imOut_temp :="1101111000000010";
when "0000000001110011"=>
    imOut_temp :="1101111000000011";
when "0000000001110100"=>
    imOut_temp :="1101111000000100";
when "0000000001110101"=>
    imOut_temp :="1101111000000101";
when "0000000001110110"=>
    imOut_temp :="1101111000000110";
when "0000000001110111"=>
    imOut_temp :="0100100000000001";
when "0000000001111000"=>
    imOut_temp :="1101111000000111";
when "0000000001111001"=>
    imOut_temp :="0100100000000001";
when "0000000001111010"=>
    imOut_temp :="1101111000001000";
when "0000000001111011"=>
    imOut_temp :="0100100000000001";
when "0000000001111100"=>
    imOut_temp :="1101111000001001";
when "0000000001111101"=>
    imOut_temp :="1110111101000000";
when "0000000001111110"=>
    imOut_temp :="0100111100000011";
when "0000000001111111"=>
    imOut_temp :="0000100000000000";
when "0000000010000000"=>
    imOut_temp :="0001000001001010";
when "0000000010000001"=>
    imOut_temp :="0110111010111111";
when "0000000010000010"=>
    imOut_temp :="0011011011000000";
when "0000000010000011"=>
    imOut_temp :="0110100001001111";
when "0000000010000100"=>
    imOut_temp :="1101111000000000";
when "0000000010000101"=>
    imOut_temp :="0000100000000000";
when "0000000010000110"=>
    imOut_temp :="1110111101000000";
when "0000000010000111"=>
    imOut_temp :="0100111100000011";
when "0000000010001000"=>
    imOut_temp :="0000100000000000";
when "0000000010001001"=>
    imOut_temp :="0001000001000001";
when "0000000010001010"=>
    imOut_temp :="0110111010111111";
when "0000000010001011"=>
    imOut_temp :="0011011011000000";
when "0000000010001100"=>
    imOut_temp :="0110100001001011";
when "0000000010001101"=>
    imOut_temp :="1101111000000000";
when "0000000010001110"=>
    imOut_temp :="0000100000000000";
when "0000000010001111"=>
    imOut_temp :="1110111101000000";
when "0000000010010000"=>
    imOut_temp :="0100111100000011";
when "0000000010010001"=>
    imOut_temp :="0000100000000000";
when "0000000010010010"=>
    imOut_temp :="0001000000111000";
when "0000000010010011"=>
    imOut_temp :="0110111010111111";
when "0000000010010100"=>
    imOut_temp :="0011011011000000";
when "0000000010010101"=>
    imOut_temp :="0110100000001010";
when "0000000010010110"=>
    imOut_temp :="1101111000000000";
when "0000000010010111"=>
    imOut_temp :="0000100000000000";
when "0000000010011000"=>
    imOut_temp :="1110111101000000";
when "0000000010011001"=>
    imOut_temp :="0100111100000011";
when "0000000010011010"=>
    imOut_temp :="0000100000000000";
when "0000000010011011"=>
    imOut_temp :="0001000000101111";
when "0000000010011100"=>
    imOut_temp :="0110111010111111";
when "0000000010011101"=>
    imOut_temp :="0011011011000000";
when "0000000010011110"=>
    imOut_temp :="0110100000001101";
when "0000000010011111"=>
    imOut_temp :="1101111000000000";
when "0000000010100000"=>
    imOut_temp :="0000100000000000";
when "0000000010100001"=>
    imOut_temp :="1110111101000000";
when "0000000010100010"=>
    imOut_temp :="0100111100000011";
when "0000000010100011"=>
    imOut_temp :="0000100000000000";
when "0000000010100100"=>
    imOut_temp :="0001000000110001";
when "0000000010100101"=>
    imOut_temp :="0000100000000000";
when "0000000010100110"=>
    imOut_temp :="0110111010111111";
when "0000000010100111"=>
    imOut_temp :="0011011011000000";
when "0000000010101000"=>
    imOut_temp :="1001111000100000";
when "0000000010101001"=>
    imOut_temp :="0110111011111111";
when "0000000010101010"=>
    imOut_temp :="1110100111001100";
when "0000000010101011"=>
    imOut_temp :="0000100000000000";
when "0000000010101100"=>
    imOut_temp :="0110100001010010";
when "0000000010101101"=>
    imOut_temp :="1110100000101010";
when "0000000010101110"=>
    imOut_temp :="0110000000110010";
when "0000000010101111"=>
    imOut_temp :="0000100000000000";
when "0000000010110000"=>
    imOut_temp :="0110100001000100";
when "0000000010110001"=>
    imOut_temp :="1110100000101010";
when "0000000010110010"=>
    imOut_temp :="0110000001001101";
when "0000000010110011"=>
    imOut_temp :="0000100000000000";
when "0000000010110100"=>
    imOut_temp :="0110100001000001";
when "0000000010110101"=>
    imOut_temp :="1110100000101010";
when "0000000010110110"=>
    imOut_temp :="0110000000001110";
when "0000000010110111"=>
    imOut_temp :="0000100000000000";
when "0000000010111000"=>
    imOut_temp :="0110100001010101";
when "0000000010111001"=>
    imOut_temp :="1110100000101010";
when "0000000010111010"=>
    imOut_temp :="0110000000000111";
when "0000000010111011"=>
    imOut_temp :="0000100000000000";
when "0000000010111100"=>
    imOut_temp :="0110100001000111";
when "0000000010111101"=>
    imOut_temp :="1110100000101010";
when "0000000010111110"=>
    imOut_temp :="0110000000001001";
when "0000000010111111"=>
    imOut_temp :="0000100000000000";
when "0000000011000000"=>
    imOut_temp :="0001011111100000";
when "0000000011000001"=>
    imOut_temp :="0000100000000000";
when "0000000011000010"=>
    imOut_temp :="0000100000000000";
when "0000000011000011"=>
    imOut_temp :="0001000011000000";
when "0000000011000100"=>
    imOut_temp :="0000100000000000";
when "0000000011000101"=>
    imOut_temp :="0000100000000000";
when "0000000011000110"=>
    imOut_temp :="0001000010000010";
when "0000000011000111"=>
    imOut_temp :="0000100000000000";
when "0000000011001000"=>
    imOut_temp :="0000100000000000";
when "0000000011001001"=>
    imOut_temp :="0001000100000011";
when "0000000011001010"=>
    imOut_temp :="0000100000000000";
when "0000000011001011"=>
    imOut_temp :="0000100000000000";
when "0000000011001100"=>
    imOut_temp :="0110111010111111";
when "0000000011001101"=>
    imOut_temp :="0011011011000000";
when "0000000011001110"=>
    imOut_temp :="0100111000000001";
when "0000000011001111"=>
    imOut_temp :="1001111000000000";
when "0000000011010000"=>
    imOut_temp :="0110111000000001";
when "0000000011010001"=>
    imOut_temp :="1110100011001100";
when "0000000011010010"=>
    imOut_temp :="0010000011111000";
when "0000000011010011"=>
    imOut_temp :="0000100000000000";
when "0000000011010100"=>
    imOut_temp :="1110111100000000";
when "0000000011010101"=>
    imOut_temp :="0000100000000000";
when "0000000011010110"=>
    imOut_temp :="0000100000000000";
when "0000000011010111"=>
    imOut_temp :="0110111010111111";
when "0000000011011000"=>
    imOut_temp :="0011011011000000";
when "0000000011011001"=>
    imOut_temp :="0100111000000001";
when "0000000011011010"=>
    imOut_temp :="1001111000000000";
when "0000000011011011"=>
    imOut_temp :="0110111000000010";
when "0000000011011100"=>
    imOut_temp :="1110100011001100";
when "0000000011011101"=>
    imOut_temp :="0010000011111000";
when "0000000011011110"=>
    imOut_temp :="0000100000000000";
when "0000000011011111"=>
    imOut_temp :="1110111100000000";
when "0000000011100000"=>
    imOut_temp :="0000100000000000";
when "0000000011100001"=>
    imOut_temp :="0110100100000110";
when "0000000011100010"=>
    imOut_temp :="0110101000000110";
when "0000000011100011"=>
    imOut_temp :="0110100010111111";
when "0000000011100100"=>
    imOut_temp :="0011000000000000";
when "0000000011100101"=>
    imOut_temp :="0100100000010000";
when "0000000011100110"=>
    imOut_temp :="1110001000101111";
when "0000000011100111"=>
    imOut_temp :="1110000001100001";
when "0000000011101000"=>
    imOut_temp :="1001100001100000";
when "0000000011101001"=>
    imOut_temp :="1110111101000000";
when "0000000011101010"=>
    imOut_temp :="0100111100000011";
when "0000000011101011"=>
    imOut_temp :="0000100000000000";
when "0000000011101100"=>
    imOut_temp :="0001011111011110";
when "0000000011101101"=>
    imOut_temp :="0000100000000000";
when "0000000011101110"=>
    imOut_temp :="0110111010111111";
when "0000000011101111"=>
    imOut_temp :="0011011011000000";
when "0000000011110000"=>
    imOut_temp :="1101111001100000";
when "0000000011110001"=>
    imOut_temp :="0011001101100011";
when "0000000011110010"=>
    imOut_temp :="1110111101000000";
when "0000000011110011"=>
    imOut_temp :="0100111100000011";
when "0000000011110100"=>
    imOut_temp :="0000100000000000";
when "0000000011110101"=>
    imOut_temp :="0001011111010101";
when "0000000011110110"=>
    imOut_temp :="0000100000000000";
when "0000000011110111"=>
    imOut_temp :="0110111010111111";
when "0000000011111000"=>
    imOut_temp :="0011011011000000";
when "0000000011111001"=>
    imOut_temp :="1101111001100000";
when "0000000011111010"=>
    imOut_temp :="0100100111111111";
when "0000000011111011"=>
    imOut_temp :="0000100000000000";
when "0000000011111100"=>
    imOut_temp :="0010100111100110";
when "0000000011111101"=>
    imOut_temp :="0000100000000000";
when "0000000011111110"=>
    imOut_temp :="0001011110100010";
when "0000000011111111"=>
    imOut_temp :="0000100000000000";
when "0000000100000000"=>
    imOut_temp :="1110111101000000";
when "0000000100000001"=>
    imOut_temp :="0100111100000011";
when "0000000100000010"=>
    imOut_temp :="0000100000000000";
when "0000000100000011"=>
    imOut_temp :="0001011111010010";
when "0000000100000100"=>
    imOut_temp :="0000100000000000";
when "0000000100000101"=>
    imOut_temp :="0110111010111111";
when "0000000100000110"=>
    imOut_temp :="0011011011000000";
when "0000000100000111"=>
    imOut_temp :="1001111010100000";
when "0000000100001000"=>
    imOut_temp :="0110111011111111";
when "0000000100001001"=>
    imOut_temp :="1110110111001100";
when "0000000100001010"=>
    imOut_temp :="0000100000000000";
when "0000000100001011"=>
    imOut_temp :="1110111101000000";
when "0000000100001100"=>
    imOut_temp :="0100111100000011";
when "0000000100001101"=>
    imOut_temp :="0000100000000000";
when "0000000100001110"=>
    imOut_temp :="0001011111000111";
when "0000000100001111"=>
    imOut_temp :="0000100000000000";
when "0000000100010000"=>
    imOut_temp :="0110111010111111";
when "0000000100010001"=>
    imOut_temp :="0011011011000000";
when "0000000100010010"=>
    imOut_temp :="1001111000100000";
when "0000000100010011"=>
    imOut_temp :="0110111011111111";
when "0000000100010100"=>
    imOut_temp :="1110100111001100";
when "0000000100010101"=>
    imOut_temp :="0000100000000000";
when "0000000100010110"=>
    imOut_temp :="0011000100100000";
when "0000000100010111"=>
    imOut_temp :="1110100110101101";
when "0000000100011000"=>
    imOut_temp :="1110111101000000";
when "0000000100011001"=>
    imOut_temp :="0100111100000011";
when "0000000100011010"=>
    imOut_temp :="0000100000000000";
when "0000000100011011"=>
    imOut_temp :="0001011110111010";
when "0000000100011100"=>
    imOut_temp :="0000100000000000";
when "0000000100011101"=>
    imOut_temp :="0110111010111111";
when "0000000100011110"=>
    imOut_temp :="0011011011000000";
when "0000000100011111"=>
    imOut_temp :="1001111010100000";
when "0000000100100000"=>
    imOut_temp :="0110111011111111";
when "0000000100100001"=>
    imOut_temp :="1110110111001100";
when "0000000100100010"=>
    imOut_temp :="0000100000000000";
when "0000000100100011"=>
    imOut_temp :="1110111101000000";
when "0000000100100100"=>
    imOut_temp :="0100111100000011";
when "0000000100100101"=>
    imOut_temp :="0000100000000000";
when "0000000100100110"=>
    imOut_temp :="0001011110101111";
when "0000000100100111"=>
    imOut_temp :="0000100000000000";
when "0000000100101000"=>
    imOut_temp :="0110111010111111";
when "0000000100101001"=>
    imOut_temp :="0011011011000000";
when "0000000100101010"=>
    imOut_temp :="1001111001000000";
when "0000000100101011"=>
    imOut_temp :="0110111011111111";
when "0000000100101100"=>
    imOut_temp :="1110101011001100";
when "0000000100101101"=>
    imOut_temp :="0000100000000000";
when "0000000100101110"=>
    imOut_temp :="0011001001000000";
when "0000000100101111"=>
    imOut_temp :="1110101010101101";
when "0000000100110000"=>
    imOut_temp :="1001100101100000";
when "0000000100110001"=>
    imOut_temp :="1110111101000000";
when "0000000100110010"=>
    imOut_temp :="0100111100000011";
when "0000000100110011"=>
    imOut_temp :="0000100000000000";
when "0000000100110100"=>
    imOut_temp :="0001011110010110";
when "0000000100110101"=>
    imOut_temp :="0000100000000000";
when "0000000100110110"=>
    imOut_temp :="0110111010111111";
when "0000000100110111"=>
    imOut_temp :="0011011011000000";
when "0000000100111000"=>
    imOut_temp :="1101111001100000";
when "0000000100111001"=>
    imOut_temp :="0011001101100011";
when "0000000100111010"=>
    imOut_temp :="1110111101000000";
when "0000000100111011"=>
    imOut_temp :="0100111100000011";
when "0000000100111100"=>
    imOut_temp :="0000100000000000";
when "0000000100111101"=>
    imOut_temp :="0001011110001101";
when "0000000100111110"=>
    imOut_temp :="0000100000000000";
when "0000000100111111"=>
    imOut_temp :="0110111010111111";
when "0000000101000000"=>
    imOut_temp :="0011011011000000";
when "0000000101000001"=>
    imOut_temp :="1101111001100000";
when "0000000101000010"=>
    imOut_temp :="0100100100000001";
when "0000000101000011"=>
    imOut_temp :="0100101011111111";
when "0000000101000100"=>
    imOut_temp :="0000100000000000";
when "0000000101000101"=>
    imOut_temp :="0010101011101010";
when "0000000101000110"=>
    imOut_temp :="0000100000000000";
when "0000000101000111"=>
    imOut_temp :="0001011101011001";
when "0000000101001000"=>
    imOut_temp :="0000100000000000";
when "0000000101001001"=>
    imOut_temp :="1110111101000000";
when "0000000101001010"=>
    imOut_temp :="0100111100000011";
when "0000000101001011"=>
    imOut_temp :="0000100000000000";
when "0000000101001100"=>
    imOut_temp :="0001011110001001";
when "0000000101001101"=>
    imOut_temp :="0000100000000000";
when "0000000101001110"=>
    imOut_temp :="0110111010111111";
when "0000000101001111"=>
    imOut_temp :="0011011011000000";
when "0000000101010000"=>
    imOut_temp :="1001111010100000";
when "0000000101010001"=>
    imOut_temp :="0110111011111111";
when "0000000101010010"=>
    imOut_temp :="1110110111001100";
when "0000000101010011"=>
    imOut_temp :="0000100000000000";
when "0000000101010100"=>
    imOut_temp :="1110111101000000";
when "0000000101010101"=>
    imOut_temp :="0100111100000011";
when "0000000101010110"=>
    imOut_temp :="0000100000000000";
when "0000000101010111"=>
    imOut_temp :="0001011101111110";
when "0000000101011000"=>
    imOut_temp :="0000100000000000";
when "0000000101011001"=>
    imOut_temp :="0110111010111111";
when "0000000101011010"=>
    imOut_temp :="0011011011000000";
when "0000000101011011"=>
    imOut_temp :="1001111000100000";
when "0000000101011100"=>
    imOut_temp :="0110111011111111";
when "0000000101011101"=>
    imOut_temp :="1110100111001100";
when "0000000101011110"=>
    imOut_temp :="0000100000000000";
when "0000000101011111"=>
    imOut_temp :="0011000100100000";
when "0000000101100000"=>
    imOut_temp :="1110100110101101";
when "0000000101100001"=>
    imOut_temp :="0110100000000000";
when "0000000101100010"=>
    imOut_temp :="1110100000101010";
when "0000000101100011"=>
    imOut_temp :="0110000000011101";
when "0000000101100100"=>
    imOut_temp :="0000100000000000";
when "0000000101100101"=>
    imOut_temp :="1110111101000000";
when "0000000101100110"=>
    imOut_temp :="0100111100000011";
when "0000000101100111"=>
    imOut_temp :="0000100000000000";
when "0000000101101000"=>
    imOut_temp :="0001011101101101";
when "0000000101101001"=>
    imOut_temp :="0000100000000000";
when "0000000101101010"=>
    imOut_temp :="0110111010111111";
when "0000000101101011"=>
    imOut_temp :="0011011011000000";
when "0000000101101100"=>
    imOut_temp :="1001111010100000";
when "0000000101101101"=>
    imOut_temp :="0110111011111111";
when "0000000101101110"=>
    imOut_temp :="1110110111001100";
when "0000000101101111"=>
    imOut_temp :="0000100000000000";
when "0000000101110000"=>
    imOut_temp :="1110111101000000";
when "0000000101110001"=>
    imOut_temp :="0100111100000011";
when "0000000101110010"=>
    imOut_temp :="0000100000000000";
when "0000000101110011"=>
    imOut_temp :="0001011101100010";
when "0000000101110100"=>
    imOut_temp :="0000100000000000";
when "0000000101110101"=>
    imOut_temp :="0110111010111111";
when "0000000101110110"=>
    imOut_temp :="0011011011000000";
when "0000000101110111"=>
    imOut_temp :="1001111001000000";
when "0000000101111000"=>
    imOut_temp :="0110111011111111";
when "0000000101111001"=>
    imOut_temp :="1110101011001100";
when "0000000101111010"=>
    imOut_temp :="0000100000000000";
when "0000000101111011"=>
    imOut_temp :="0011001001000000";
when "0000000101111100"=>
    imOut_temp :="1110101010101101";
when "0000000101111101"=>
    imOut_temp :="1101100101000000";
when "0000000101111110"=>
    imOut_temp :="0000100000000000";
when "0000000101111111"=>
    imOut_temp :="0001011111001001";
when "0000000110000000"=>
    imOut_temp :="0000100000000000";
when "0000000110000001"=>
    imOut_temp :="0000100000000000";
when "0000000110000010"=>
    imOut_temp :="0001011100011110";
when "0000000110000011"=>
    imOut_temp :="0000100000000000";
when "0000000110000100"=>
    imOut_temp :="1110111101000000";
when "0000000110000101"=>
    imOut_temp :="0100111100000011";
when "0000000110000110"=>
    imOut_temp :="0000100000000000";
when "0000000110000111"=>
    imOut_temp :="0001011101001110";
when "0000000110001000"=>
    imOut_temp :="0000100000000000";
when "0000000110001001"=>
    imOut_temp :="0110111010111111";
when "0000000110001010"=>
    imOut_temp :="0011011011000000";
when "0000000110001011"=>
    imOut_temp :="1001111010100000";
when "0000000110001100"=>
    imOut_temp :="0110111011111111";
when "0000000110001101"=>
    imOut_temp :="1110110111001100";
when "0000000110001110"=>
    imOut_temp :="0000100000000000";
when "0000000110001111"=>
    imOut_temp :="1110111101000000";
when "0000000110010000"=>
    imOut_temp :="0100111100000011";
when "0000000110010001"=>
    imOut_temp :="0000100000000000";
when "0000000110010010"=>
    imOut_temp :="0001011101000011";
when "0000000110010011"=>
    imOut_temp :="0000100000000000";
when "0000000110010100"=>
    imOut_temp :="0110111010111111";
when "0000000110010101"=>
    imOut_temp :="0011011011000000";
when "0000000110010110"=>
    imOut_temp :="1001111000100000";
when "0000000110010111"=>
    imOut_temp :="0110111011111111";
when "0000000110011000"=>
    imOut_temp :="1110100111001100";
when "0000000110011001"=>
    imOut_temp :="0000100000000000";
when "0000000110011010"=>
    imOut_temp :="0011000100100000";
when "0000000110011011"=>
    imOut_temp :="1110100110101101";
when "0000000110011100"=>
    imOut_temp :="1110111101000000";
when "0000000110011101"=>
    imOut_temp :="0100111100000011";
when "0000000110011110"=>
    imOut_temp :="0000100000000000";
when "0000000110011111"=>
    imOut_temp :="0001011100110110";
when "0000000110100000"=>
    imOut_temp :="0000100000000000";
when "0000000110100001"=>
    imOut_temp :="0110111010111111";
when "0000000110100010"=>
    imOut_temp :="0011011011000000";
when "0000000110100011"=>
    imOut_temp :="1001111010100000";
when "0000000110100100"=>
    imOut_temp :="0110111011111111";
when "0000000110100101"=>
    imOut_temp :="1110110111001100";
when "0000000110100110"=>
    imOut_temp :="0000100000000000";
when "0000000110100111"=>
    imOut_temp :="1110111101000000";
when "0000000110101000"=>
    imOut_temp :="0100111100000011";
when "0000000110101001"=>
    imOut_temp :="0000100000000000";
when "0000000110101010"=>
    imOut_temp :="0001011100101011";
when "0000000110101011"=>
    imOut_temp :="0000100000000000";
when "0000000110101100"=>
    imOut_temp :="0110111010111111";
when "0000000110101101"=>
    imOut_temp :="0011011011000000";
when "0000000110101110"=>
    imOut_temp :="1001111001000000";
when "0000000110101111"=>
    imOut_temp :="0110111011111111";
when "0000000110110000"=>
    imOut_temp :="1110101011001100";
when "0000000110110001"=>
    imOut_temp :="0000100000000000";
when "0000000110110010"=>
    imOut_temp :="0011001001000000";
when "0000000110110011"=>
    imOut_temp :="1110101010101101";
when "0000000110110100"=>
    imOut_temp :="1001100101100000";
when "0000000110110101"=>
    imOut_temp :="1110111101000000";
when "0000000110110110"=>
    imOut_temp :="0100111100000011";
when "0000000110110111"=>
    imOut_temp :="0000100000000000";
when "0000000110111000"=>
    imOut_temp :="0001011100010010";
when "0000000110111001"=>
    imOut_temp :="0000100000000000";
when "0000000110111010"=>
    imOut_temp :="0110111010111111";
when "0000000110111011"=>
    imOut_temp :="0011011011000000";
when "0000000110111100"=>
    imOut_temp :="1101111001100000";
when "0000000110111101"=>
    imOut_temp :="0011001101100011";
when "0000000110111110"=>
    imOut_temp :="1110111101000000";
when "0000000110111111"=>
    imOut_temp :="0100111100000011";
when "0000000111000000"=>
    imOut_temp :="0000100000000000";
when "0000000111000001"=>
    imOut_temp :="0001011100001001";
when "0000000111000010"=>
    imOut_temp :="0000100000000000";
when "0000000111000011"=>
    imOut_temp :="0110111010111111";
when "0000000111000100"=>
    imOut_temp :="0011011011000000";
when "0000000111000101"=>
    imOut_temp :="1101111001100000";
when "0000000111000110"=>
    imOut_temp :="0100100100000001";
when "0000000111000111"=>
    imOut_temp :="0100101011111111";
when "0000000111001000"=>
    imOut_temp :="0000100000000000";
when "0000000111001001"=>
    imOut_temp :="0010101011101010";
when "0000000111001010"=>
    imOut_temp :="0000100000000000";
when "0000000111001011"=>
    imOut_temp :="0001011011010101";
when "0000000111001100"=>
    imOut_temp :="0000100000000000";
when "0000000111001101"=>
    imOut_temp :="1110111101000000";
when "0000000111001110"=>
    imOut_temp :="0100111100000011";
when "0000000111001111"=>
    imOut_temp :="0000100000000000";
when "0000000111010000"=>
    imOut_temp :="0001011100000101";
when "0000000111010001"=>
    imOut_temp :="0000100000000000";
when "0000000111010010"=>
    imOut_temp :="0110111010111111";
when "0000000111010011"=>
    imOut_temp :="0011011011000000";
when "0000000111010100"=>
    imOut_temp :="1001111010100000";
when "0000000111010101"=>
    imOut_temp :="0110111011111111";
when "0000000111010110"=>
    imOut_temp :="1110110111001100";
when "0000000111010111"=>
    imOut_temp :="0000100000000000";
when "0000000111011000"=>
    imOut_temp :="1110111101000000";
when "0000000111011001"=>
    imOut_temp :="0100111100000011";
when "0000000111011010"=>
    imOut_temp :="0000100000000000";
when "0000000111011011"=>
    imOut_temp :="0001011011111010";
when "0000000111011100"=>
    imOut_temp :="0000100000000000";
when "0000000111011101"=>
    imOut_temp :="0110111010111111";
when "0000000111011110"=>
    imOut_temp :="0011011011000000";
when "0000000111011111"=>
    imOut_temp :="1001111001000000";
when "0000000111100000"=>
    imOut_temp :="0110111011111111";
when "0000000111100001"=>
    imOut_temp :="1110101011001100";
when "0000000111100010"=>
    imOut_temp :="0000100000000000";
when "0000000111100011"=>
    imOut_temp :="0011001001000000";
when "0000000111100100"=>
    imOut_temp :="1110101010101101";
when "0000000111100101"=>
    imOut_temp :="0100001011000000";
when "0000000111100110"=>
    imOut_temp :="0110111110111111";
when "0000000111100111"=>
    imOut_temp :="0011011111100000";
when "0000000111101000"=>
    imOut_temp :="0100111100010000";
when "0000000111101001"=>
    imOut_temp :="1001111110100101";
when "0000000111101010"=>
    imOut_temp :="0110001111111111";
when "0000000111101011"=>
    imOut_temp :="1101010100000000";
when "0000000111101100"=>
    imOut_temp :="1111010100000000";
when "0000000111101101"=>
    imOut_temp :="0110100110000000";
when "0000000111101110"=>
    imOut_temp :="0011000100100000";
when "0000000111101111"=>
    imOut_temp :="1110110100101101";
when "0000000111110000"=>
    imOut_temp :="1001111100000000";
when "0000000111110001"=>
    imOut_temp :="1001111100100001";
when "0000000111110010"=>
    imOut_temp :="1001111101000010";
when "0000000111110011"=>
    imOut_temp :="1001111101100011";
when "0000000111110100"=>
    imOut_temp :="1001111110000100";
when "0000000111110101"=>
    imOut_temp :="1110111101000000";
when "0000000111110110"=>
    imOut_temp :="0100111100000100";
when "0000000111110111"=>
    imOut_temp :="1111010100000001";
when "0000000111111000"=>
    imOut_temp :="1110111000000000";
when "0000000111111001"=>
    imOut_temp :="1001010100000000";
when "0000000111111010"=>
    imOut_temp :="0000100000000000";
when "0000000111111011"=>
    imOut_temp :="0000100000000000";
when "0000000111111100"=>
    imOut_temp :="0110001100000001";
when "0000000111111101"=>
    imOut_temp :="0110111110111111";
when "0000000111111110"=>
    imOut_temp :="0011011111100000";
when "0000000111111111"=>
    imOut_temp :="0100111100010000";
when "0000001000000000"=>
    imOut_temp :="1101111100000000";
when "0000001000000001"=>
    imOut_temp :="1101111100100001";
when "0000001000000010"=>
    imOut_temp :="1101111101000010";
when "0000001000000011"=>
    imOut_temp :="1101111101100011";
when "0000001000000100"=>
    imOut_temp :="1101111110000100";
when "0000001000000101"=>
    imOut_temp :="1101111110100101";
when "0000001000000110"=>
    imOut_temp :="1111000000000000";
when "0000001000000111"=>
    imOut_temp :="0110100101111111";
when "0000001000001000"=>
    imOut_temp :="0011000100100000";
when "0000001000001001"=>
    imOut_temp :="0110101011111111";
when "0000001000001010"=>
    imOut_temp :="1110100101001101";
when "0000001000001011"=>
    imOut_temp :="1110100000101100";
when "0000001000001100"=>
    imOut_temp :="1111000000000001";
when "0000001000001101"=>
    imOut_temp :="0110100100000111";
when "0000001000001110"=>
    imOut_temp :="1110111101000000";
when "0000001000001111"=>
    imOut_temp :="0100111100000011";
when "0000001000010000"=>
    imOut_temp :="0000100000000000";
when "0000001000010001"=>
    imOut_temp :="0001011010111001";
when "0000001000010010"=>
    imOut_temp :="0000100000000000";
when "0000001000010011"=>
    imOut_temp :="0110111010111111";
when "0000001000010100"=>
    imOut_temp :="0011011011000000";
when "0000001000010101"=>
    imOut_temp :="1101111000100000";
when "0000001000010110"=>
    imOut_temp :="0001011010001010";
when "0000001000010111"=>
    imOut_temp :="0000100000000000";
----chuankou
--when "1011111100000000"=>
--	imOut_temp := "0000000000000001";
--when "1011111100000001"=>
--	imOut_temp := "0000000000000001";
--					when "0000000000000000"=>
--						imOut_temp := "0110100000100000";
--					when "0000000000000001"=>
--						imOut_temp := "1101100000000000";
--					when "0000000000000010"=>
--						imOut_temp := "1101100000000001";
--					when "0000000000000011"=>
--						imOut_temp := "1101100000000010";
--					when "0000000000000100"=>
--						imOut_temp := "1101100000000011";
--					when "0000000000000101"=>
--						imOut_temp := "1101100000000100";
--					when "0000000000000110"=>
--						imOut_temp := "1101100000000101";
--					when "0000000000000111"=>
--						imOut_temp := "1101100000000110";
--					when "0000000000001000"=>
--						imOut_temp := "0100100100000001";
--					when "0000000000001001"=>
--						imOut_temp := "1101100000100111";
--					when "0000000000001010"=>
--						imOut_temp := "0100100100000001";
--					when "0000000000001011"=>
--						imOut_temp := "1101100000101000";
					when others=>
						imOut_temp := "0000100000000000";
				end case;
				end if;
			end if;
			
		end if;
	end process;
	process(clk,rst)
	begin
		if(rst = '0') then
			dmOut <= "0000000000000000";
			ImOut <= "0000100000000000";
			req_stall_im <= '0';
			--req_stall_dm <= '0';
			--display_im <= "0000000000000000";
			--display_dm <= "0000000000000000";
		elsif(falling_edge(clk)) then
			req_stall_im <= '0';
			--req_stall_dm <= '0';
			imOut <= imOut_temp;
			if(state_keep = '1') then
				dmOut <= (others=>'1');
			else
				dmOut <= dmOut_temp;
			 
			end if;
		end if;
	end process;
end Behavioral;

